module cnt_6();
input rst, clk;
output q;
reg temp;

always@(negedge rst, posedge clk) begin


end

endmodule
