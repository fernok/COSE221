module MUX(A, B, C, D, s, out);
input [4:0] A, B, C, D;
input [1:0] s;
output reg [4:0] out;

always@(s, A, B, C, D)
begin
case(s)
	2'b00 : out = A;
	2'b01 : out = B;
	2'b10 : out = C;
	2'b11 : out = D;
endcase
end

endmodule
