module cnt24(rst, in_clk, h1, h10);
input rst, in_clk;
output reg [3:0] h1, h10;
reg [4:0] q, temp;

always@(negedge rst, posedge in_clk)
begin
if(!rst)
   begin
      q <= 0;
      temp <= 0;
   end
else
   begin
      if(temp == 23)
         temp <= 0;
      else
         temp <= temp + 1;
      q <= temp;
   end
end

always@(q)
begin
if(q < 10)
   begin
      h10 <= 0;
      h1 <= q;
   end
else if(10 <= q && q < 20)
   begin
      h10 <= 1;
      h1 <= q - 10;
   end
else if(20 <= q)
   begin
      h10 <= 2;
      h1 <= q - 20;
   end
end
endmodule
