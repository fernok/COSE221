module Fourbit(A, B, EQ, ALB, AGB);
input [3:0] A, B;
output reg EQ, ALB, AGB;
wire [3:0] x;

assign x[0] = (A[0]&B[0])|(~A[0]*~B[0]);
assign x[1] = (A[1]&B[1])|(~A[1]*~B[1]);
assign x[2] = (A[2]&B[2])|(~A[2]*~B[2]);
assign x[3] = (A[3]&B[3])|(~A[3]*~B[3]);

always@(A, B, x)
begin
if(x[3]&x[2]&x[1]&x[0]) 
begin EQ = 1; ALB = 0; AGB = 0; end 
else if((A[3]&~B[3])|(x[3]&A[2]&~B[2])|(x[3]&x[2]&A[1]&~B[1])|(x[3]&x[2]&x[1]&A[0]&~B[0]))
begin EQ = 0; ALB = 0; AGB = 1; end
else 
begin EQ = 0; ALB = 1; AGB = 0; end
end

endmodule
